library ieee;

use ieee.numeric_std.all;
use work.cpu_defs_pack.all;
use work.bit_vector_natural_pack.all;

entity srli_s is
    port(
        a: in datatype; --data form rs1
        b: in datatype; --zero extended lower five bit of rs2 (shamt)
        c: out datatype --data in rd
    );

end entity;

architecture behav of srli_s is
    signal shift: integer;

    begin
        
        shift <= bit_vector2natural(b);

        process(a, b)
            variable temp: datatype;
        begin
    
            if (shift > 31) then
                c <= (others => '0');
                
            else
                for i in 1 to shift loop
                    temp := '0' & a(datasize-1 downto 1);
                end loop;
                --c <= (others => '0') & a[31 downt shift];
        	c <= temp;
            end if;
		
        end process;
	
end architecture;